`timescale 	1ns				/ 100ps

`include "demux_estructural.v"
`include "demux_conductual.v"
`include "probador.v"

module banco_pruebas_conductual; // Testbench

    wire [3:0] data_out0_ESTRUC, data_out1_ESTRUC, data_out0_COND,data_out1_COND,data_in;
	wire clk, reset_L;

	demux_conductual	demux_conduct(	/*AUTOINST*/
					      // Outputs
					      .data_out0	(data_out0_COND[3:0]),
					      .data_out1	(data_out1_COND[3:0]),
					      // Inputs
					      .clk		(clk),
					      .reset_L		(reset_L),
					      .data_in		(data_in[3:0]));

	// Descripci�n conductual de alarma
	demux_estructural	demux_estruc(	/*AUTOINST*/
					     // Outputs
					     .data_out0		(data_out0_ESTRUC[3:0]),
					     .data_out1		(data_out1_ESTRUC[3:0]),
					     // Inputs
					     .clk		(clk),
					     .reset_L		(reset_L),
					     .data_in		(data_in[3:0]));

	// Probador: generador de se�ales y monitor
	probador probador_(     /*AUTOINST*/
			   // Outputs
			   .data_in		(data_in[3:0]),
			   .reset_L		(reset_L),
			   .clk			(clk),
			   // Inputs
			   .data_out0_ESTRUC	(data_out0_ESTRUC[3:0]),
			   .data_out1_ESTRUC	(data_out1_ESTRUC[3:0]),
			   .data_out0_COND	(data_out0_COND[3:0]),
			   .data_out1_COND	(data_out1_COND[3:0]));
endmodule
