//Generador de señales y monitor de datos
module probador( 
	output reg	[7:0]			data_in_0,
	output reg 					valid_in_0,
	output reg	[7:0]			data_in_1,
	output reg 					valid_in_1,
	output reg 					reset,	
	output reg 					clk8f,
	input 		[7:0]			data_out_0_c,
	input 	 					valid_out_0_c,
	input 		[7:0]			data_out_1_c,
	input 	 					valid_out_1_c,
	input 		[7:0]			data_out_0_s,
	input 	 					valid_out_0_s,
	input 		[7:0]			data_out_1_s,
	input 	 					valid_out_1_s,
	input						clk4f,
	input						clk2f,
	input						clkf);

	
	initial begin
		$dumpfile("proy1.vcd"); //Archivo de dump
		$dumpvars;				//Ordena dumpear variables a demux.vcd
		
		$display ("\t\t\tclk,\tclks,\treset");	//Mensaje inicial que se imprime en consola
		
		$monitor($time,"\t%b\t%b\t\t%b\t\t%b\t%b", clk8f, clkf, clk2f, clk4f, reset); //Valores que se imprimen con cada cambio 

		data_in_0 = 0;		//A continuaci�n, se generan las se�ales de prueba a usar para la simulaci�n	
		data_in_1 = 0;
		valid_in_0 = 0;
		valid_in_1 = 0;
		reset = 0;
		@(posedge clk8f);
		data_in_0 <= 'h11;
		data_in_1 <= 'hFF;
		@(posedge clk8f);
		data_in_0 <= 'h11;
		data_in_1 <= 'hFF;
		@(posedge clk8f);
		data_in_0 <= 'h11;
		data_in_1 <= 'hFF;
		@(posedge clk8f);
		data_in_0 <= 'h11;
		data_in_1 <= 'hFF;
		reset <= 1;
		@(posedge clk8f);
		data_in_0 <= 'h12;
		data_in_1 <= 'hFE;
		@(posedge clk8f);
		data_in_0 <= 'h12;
		data_in_1 <= 'hFE;
		@(posedge clk8f);
		data_in_0 <= 'h12;
		data_in_1 <= 'hFE;
		@(posedge clk8f);
		data_in_0 <= 'h12;
		data_in_1 <= 'hFE;
		@(posedge clk8f);
		data_in_0 <= 'h12;
		data_in_1 <= 'hFE;
		@(posedge clk8f);
		data_in_0 <= 'h12;
		data_in_1 <= 'hFE;
		@(posedge clk8f);
		data_in_0 <= 'h12;
		data_in_1 <= 'hFE;
		@(posedge clk8f);
		data_in_0 <= 'h12;
		data_in_1 <= 'hFE;
		@(posedge clk8f);
		data_in_0 <= 'h13;
		data_in_1 <= 'hFD;
		valid_in_0 <= 1;
		@(posedge clk8f);
		data_in_0 <= 'h13;
		data_in_1 <= 'hFD;
		valid_in_0 <= 1;
		@(posedge clk8f);
		data_in_0 <= 'h13;
		data_in_1 <= 'hFD;
		valid_in_0 <= 1;
		@(posedge clk8f);
		data_in_0 <= 'h13;
		data_in_1 <= 'hFD;		
		valid_in_0 <= 1;
		@(posedge clk8f);
		data_in_0 <= 'h13;
		data_in_1 <= 'hFD;
		valid_in_0 <= 1;
		@(posedge clk8f);
		data_in_0 <= 'h13;
		data_in_1 <= 'hFD;
		valid_in_0 <= 1;
		@(posedge clk8f);
		data_in_0 <= 'h13;
		data_in_1 <= 'hFD;
		valid_in_0 <= 1;
		@(posedge clk8f);
		data_in_0 <= 'h13;
		data_in_1 <= 'hFD;		
		valid_in_0 <= 1;
		@(posedge clk8f);
		data_in_0 <= 'h14;
		data_in_1 <= 'hFC;
		@(posedge clk8f);
		data_in_0 <= 'h14;
		data_in_1 <= 'hFC;
		@(posedge clk8f);
		data_in_0 <= 'h14;
		data_in_1 <= 'hFC;
		@(posedge clk8f);
		data_in_0 <= 'h14;
		data_in_1 <= 'hFC;
		@(posedge clk8f);
		data_in_0 <= 'h14;
		data_in_1 <= 'hFC;
		@(posedge clk8f);
		data_in_0 <= 'h14;
		data_in_1 <= 'hFC;
		@(posedge clk8f);
		data_in_0 <= 'h14;
		data_in_1 <= 'hFC;
		@(posedge clk8f);
		data_in_0 <= 'h14;
		data_in_1 <= 'hFC;
		@(posedge clk8f);
		data_in_0 <= 'h15;
		data_in_1 <= 'hFB;
		valid_in_0 <= 0;
		@(posedge clk8f);
		data_in_0 <= 'h15;
		data_in_1 <= 'hFB;
		valid_in_0 <= 0;
		@(posedge clk8f);
		data_in_0 <= 'h15;
		data_in_1 <= 'hFB;
		valid_in_0 <= 0;
		@(posedge clk8f);
		data_in_0 <= 'h15;
		data_in_1 <= 'hFB;
		valid_in_0 <= 0;
		@(posedge clk8f);
		data_in_0 <= 'h15;
		data_in_1 <= 'hFB;
		valid_in_0 <= 0;
		@(posedge clk8f);
		data_in_0 <= 'h15;
		data_in_1 <= 'hFB;
		valid_in_0 <= 0;
		@(posedge clk8f);
		data_in_0 <= 'h15;
		data_in_1 <= 'hFB;
		valid_in_0 <= 0;
		@(posedge clk8f);
		data_in_0 <= 'h15;
		data_in_1 <= 'hFB;
		valid_in_0 <= 0;
		@(posedge clk8f);
		data_in_0 <= 'h16;
		data_in_1 <= 'hFA;
		@(posedge clk8f);
		data_in_0 <= 'h16;
		data_in_1 <= 'hFA;
		@(posedge clk8f);
		data_in_0 <= 'h16;
		data_in_1 <= 'hFA;
		@(posedge clk8f);
		data_in_0 <= 'h16;
		data_in_1 <= 'hFA;
		@(posedge clk8f);
		data_in_0 <= 'h16;
		data_in_1 <= 'hFA;
		@(posedge clk8f);
		data_in_0 <= 'h16;
		data_in_1 <= 'hFA;
		@(posedge clk8f);
		data_in_0 <= 'h16;
		data_in_1 <= 'hFA;
		@(posedge clk8f);
		data_in_0 <= 'h16;
		data_in_1 <= 'hFA;
		@(posedge clk8f);
		data_in_0 <= 'h17;
		data_in_1 <= 'hF9;
		valid_in_1 <= 1;
		@(posedge clk8f);
		data_in_0 <= 'h17;
		data_in_1 <= 'hF9;
		valid_in_1 <= 1;
		@(posedge clk8f);
		data_in_0 <= 'h17;
		data_in_1 <= 'hF9;
		valid_in_1 <= 1;
		@(posedge clk8f);
		data_in_0 <= 'h17;
		data_in_1 <= 'hF9;
		valid_in_1 <= 1;
		@(posedge clk8f);
		data_in_0 <= 'h17;
		data_in_1 <= 'hF9;
		valid_in_1 <= 1;
		@(posedge clk8f);
		data_in_0 <= 'h17;
		data_in_1 <= 'hF9;
		valid_in_1 <= 1;
		@(posedge clk8f);
		data_in_0 <= 'h17;
		data_in_1 <= 'hF9;
		valid_in_1 <= 1;
		@(posedge clk8f);
		data_in_0 <= 'h17;
		data_in_1 <= 'hF9;
		valid_in_1 <= 1;
		@(posedge clk8f);
		data_in_0 <= 'h18;
		data_in_1 <= 'hF8;
		@(posedge clk8f);
		data_in_0 <= 'h18;
		data_in_1 <= 'hF8;
		@(posedge clk8f);
		data_in_0 <= 'h18;
		data_in_1 <= 'hF8;
		@(posedge clk8f);
		data_in_0 <= 'h18;
		data_in_1 <= 'hF8;
		@(posedge clk8f);
		data_in_0 <= 'h18;
		data_in_1 <= 'hF8;
		@(posedge clk8f);
		data_in_0 <= 'h18;
		data_in_1 <= 'hF8;
		@(posedge clk8f);
		data_in_0 <= 'h18;
		data_in_1 <= 'hF8;
		@(posedge clk8f);
		data_in_0 <= 'h18;
		data_in_1 <= 'hF8;
		@(posedge clk8f);
		data_in_0 <= 'h19;
		data_in_1 <= 'hF7;
		valid_in_1 <= 0;
		@(posedge clk8f);
		data_in_0 <= 'h19;
		data_in_1 <= 'hF7;
		valid_in_1 <= 0;
		@(posedge clk8f);
		data_in_0 <= 'h19;
		data_in_1 <= 'hF7;
		valid_in_1 <= 0;
		@(posedge clk8f);
		data_in_0 <= 'h19;
		data_in_1 <= 'hF7;
		valid_in_1 <= 0;
		@(posedge clk8f);
		data_in_0 <= 'h19;
		data_in_1 <= 'hF7;
		valid_in_1 <= 0;
		@(posedge clk8f);
		data_in_0 <= 'h19;
		data_in_1 <= 'hF7;
		valid_in_1 <= 0;
		@(posedge clk8f);
		data_in_0 <= 'h19;
		data_in_1 <= 'hF7;
		valid_in_1 <= 0;
		@(posedge clk8f);
		data_in_0 <= 'h19;
		data_in_1 <= 'hF7;
		valid_in_1 <= 0;
		@(posedge clk8f);
		data_in_0 <= 'h1A;
		data_in_1 <= 'hF6;
		@(posedge clk8f);
		data_in_0 <= 'h1A;
		data_in_1 <= 'hF6;
		@(posedge clk8f);
		data_in_0 <= 'h1A;
		data_in_1 <= 'hF6;
		@(posedge clk8f);
		data_in_0 <= 'h1A;
		data_in_1 <= 'hF6;
		@(posedge clk8f);
		data_in_0 <= 'h1A;
		data_in_1 <= 'hF6;
		@(posedge clk8f);
		data_in_0 <= 'h1A;
		data_in_1 <= 'hF6;
		@(posedge clk8f);
		data_in_0 <= 'h1A;
		data_in_1 <= 'hF6;
		@(posedge clk8f);
		data_in_0 <= 'h1A;
		data_in_1 <= 'hF6;
		@(posedge clk8f);
		data_in_0 <= 'h1B;
		data_in_1 <= 'hF5;
		valid_in_0 <= 1;		
		valid_in_1 <= 1;
		@(posedge clk8f);
		data_in_0 <= 'h1B;
		data_in_1 <= 'hF5;
		@(posedge clk8f);
		data_in_0 <= 'h1B;
		data_in_1 <= 'hF5;
		@(posedge clk8f);
		data_in_0 <= 'h1B;
		data_in_1 <= 'hF5;
		@(posedge clk8f);
		data_in_0 <= 'h1B;
		data_in_1 <= 'hF5;
		@(posedge clk8f);
		data_in_0 <= 'h1B;
		data_in_1 <= 'hF5;
		@(posedge clk8f);
		data_in_0 <= 'h1B;
		data_in_1 <= 'hF5;
		@(posedge clk8f);
		data_in_0 <= 'h1B;
		data_in_1 <= 'hF5;
		@(posedge clk8f);
		data_in_0 <= 'h1C;
		data_in_1 <= 'hF4;		
		valid_in_1 <= 0;
		@(posedge clk8f);
		data_in_0 <= 'h1C;
		data_in_1 <= 'hF4;
		@(posedge clk8f);
		data_in_0 <= 'h1C;
		data_in_1 <= 'hF4;
		@(posedge clk8f);
		data_in_0 <= 'h1C;
		data_in_1 <= 'hF4;
		@(posedge clk8f);
		data_in_0 <= 'h1C;
		data_in_1 <= 'hF4;
		@(posedge clk8f);
		data_in_0 <= 'h1C;
		data_in_1 <= 'hF4;
		@(posedge clk8f);
		data_in_0 <= 'h1C;
		data_in_1 <= 'hF4;
		@(posedge clk8f);
		data_in_0 <= 'h1C;
		data_in_1 <= 'hF4;
		@(posedge clk8f);
		data_in_0 <= 'h1D;
		data_in_1 <= 'hF3;
		valid_in_0 <= 0;
		@(posedge clk8f);
		data_in_0 <= 'h1D;
		data_in_1 <= 'hF3;
		@(posedge clk8f);
		data_in_0 <= 'h1D;
		data_in_1 <= 'hF3;
		@(posedge clk8f);
		data_in_0 <= 'h1D;
		data_in_1 <= 'hF3;
		@(posedge clk8f);
		data_in_0 <= 'h1D;
		data_in_1 <= 'hF3;
		@(posedge clk8f);
		data_in_0 <= 'h1D;
		data_in_1 <= 'hF3;
		@(posedge clk8f);
		data_in_0 <= 'h1D;
		data_in_1 <= 'hF3;
		@(posedge clk8f);
		data_in_0 <= 'h1D;
		data_in_1 <= 'hF3;
		@(posedge clk8f);
		data_in_0 <= 'h1E;
		data_in_1 <= 'hF2;
		@(posedge clk8f);
		data_in_0 <= 'h1E;
		data_in_1 <= 'hF2;
		@(posedge clk8f);
		data_in_0 <= 'h1E;
		data_in_1 <= 'hF2;
		@(posedge clk8f);
		data_in_0 <= 'h1E;
		data_in_1 <= 'hF2;
		@(posedge clk8f);
		data_in_0 <= 'h1E;
		data_in_1 <= 'hF2;
		@(posedge clk8f);
		data_in_0 <= 'h1E;
		data_in_1 <= 'hF2;
		@(posedge clk8f);
		data_in_0 <= 'h1E;
		data_in_1 <= 'hF2;
		@(posedge clk8f);
		data_in_0 <= 'h1E;
		data_in_1 <= 'hF2;
		@(posedge clk8f);
		data_in_0 <= 'h1F;
		data_in_1 <= 'hF1;
		valid_in_0 <= 1;
		valid_in_1 <= 1;
		@(posedge clk8f);
		data_in_0 <= 'h1F;
		data_in_1 <= 'hF1;
		@(posedge clk8f);
		data_in_0 <= 'h1F;
		data_in_1 <= 'hF1;
		@(posedge clk8f);
		data_in_0 <= 'h1F;
		data_in_1 <= 'hF1;
		@(posedge clk8f);
		data_in_0 <= 'h1F;
		data_in_1 <= 'hF1;
		@(posedge clk8f);
		data_in_0 <= 'h1F;
		data_in_1 <= 'hF1;
		@(posedge clk8f);
		data_in_0 <= 'h1F;
		data_in_1 <= 'hF1;
		@(posedge clk8f);
		data_in_0 <= 'h1F;
		data_in_1 <= 'hF1;
		@(posedge clk8f);
		data_in_0 <= 'h20;
		data_in_1 <= 'hF0;
		valid_in_1 <= 0;
		@(posedge clk8f);
		data_in_0 <= 'h20;
		data_in_1 <= 'hF0;
		@(posedge clk8f);
		data_in_0 <= 'h20;
		data_in_1 <= 'hF0;
		@(posedge clk8f);
		data_in_0 <= 'h20;
		data_in_1 <= 'hF0;
		@(posedge clk8f);
		data_in_0 <= 'h20;
		data_in_1 <= 'hF0;
		@(posedge clk8f);
		data_in_0 <= 'h20;
		data_in_1 <= 'hF0;
		@(posedge clk8f);
		data_in_0 <= 'h20;
		data_in_1 <= 'hF0;
		@(posedge clk8f);
		data_in_0 <= 'h20;
		data_in_1 <= 'hF0;
		@(posedge clk8f);
		data_in_0 <= 'h21;
		data_in_1 <= 'hEF;
		valid_in_0 <= 0;
		@(posedge clk8f);
		data_in_0 <= 'h21;
		data_in_1 <= 'hEF;
		@(posedge clk8f);
		data_in_0 <= 'h21;
		data_in_1 <= 'hEF;
		@(posedge clk8f);
		data_in_0 <= 'h21;
		data_in_1 <= 'hEF;
		@(posedge clk8f);
		data_in_0 <= 'h21;
		data_in_1 <= 'hEF;
		@(posedge clk8f);
		data_in_0 <= 'h21;
		data_in_1 <= 'hEF;
		@(posedge clk8f);
		data_in_0 <= 'h21;
		data_in_1 <= 'hEF;
		@(posedge clk8f);
		data_in_0 <= 'h21;
		data_in_1 <= 'hEF;
		@(posedge clk8f);
		data_in_0 <= 'h22;
		data_in_1 <= 'hEE;
		@(posedge clk8f);
		data_in_0 <= 'h22;
		data_in_1 <= 'hEE;
		@(posedge clk8f);
		data_in_0 <= 'h22;
		data_in_1 <= 'hEE;
		@(posedge clk8f);
		data_in_0 <= 'h22;
		data_in_1 <= 'hEE;
		@(posedge clk8f);
		data_in_0 <= 'h22;
		data_in_1 <= 'hEE;
		@(posedge clk8f);
		data_in_0 <= 'h22;
		data_in_1 <= 'hEE;
		@(posedge clk8f);
		data_in_0 <= 'h22;
		data_in_1 <= 'hEE;
		@(posedge clk8f);
		data_in_0 <= 'h22;
		data_in_1 <= 'hEE;
		@(posedge clk8f);
		data_in_0 <= 'h23;
		data_in_1 <= 'hED;
		valid_in_0 <= 1;
		valid_in_1 <= 1;
		@(posedge clk8f);
		data_in_0 <= 'h23;
		data_in_1 <= 'hED;
		@(posedge clk8f);
		data_in_0 <= 'h23;
		data_in_1 <= 'hED;
		@(posedge clk8f);
		data_in_0 <= 'h23;
		data_in_1 <= 'hED;
		@(posedge clk8f);
		data_in_0 <= 'h23;
		data_in_1 <= 'hED;
		@(posedge clk8f);
		data_in_0 <= 'h23;
		data_in_1 <= 'hED;
		@(posedge clk8f);
		data_in_0 <= 'h23;
		data_in_1 <= 'hED;
		@(posedge clk8f);
		data_in_0 <= 'h23;
		data_in_1 <= 'hED;
		@(posedge clk8f);
		data_in_0 <= 'h24;
		data_in_1 <= 'hEC;
		valid_in_0 <= 0;
		@(posedge clk8f);
		data_in_0 <= 'h24;
		data_in_1 <= 'hEC;
		@(posedge clk8f);
		data_in_0 <= 'h24;
		data_in_1 <= 'hEC;
		@(posedge clk8f);
		data_in_0 <= 'h24;
		data_in_1 <= 'hEC;
		@(posedge clk8f);
		data_in_0 <= 'h24;
		data_in_1 <= 'hEC;
		@(posedge clk8f);
		data_in_0 <= 'h24;
		data_in_1 <= 'hEC;
		@(posedge clk8f);
		data_in_0 <= 'h24;
		data_in_1 <= 'hEC;
		@(posedge clk8f);
		data_in_0 <= 'h24;
		data_in_1 <= 'hEC;
		@(posedge clk8f);
		data_in_0 <= 'h25;
		data_in_1 <= 'hEB;
		valid_in_1 <= 0;
		@(posedge clk8f);
		data_in_0 <= 'h25;
		data_in_1 <= 'hEB;
		@(posedge clk8f);
		data_in_0 <= 'h25;
		data_in_1 <= 'hEB;
		@(posedge clk8f);
		data_in_0 <= 'h25;
		data_in_1 <= 'hEB;
		@(posedge clk8f);
		data_in_0 <= 'h25;
		data_in_1 <= 'hEB;
		@(posedge clk8f);
		data_in_0 <= 'h25;
		data_in_1 <= 'hEB;
		@(posedge clk8f);
		data_in_0 <= 'h25;
		data_in_1 <= 'hEB;
		@(posedge clk8f);
		data_in_0 <= 'h25;
		data_in_1 <= 'hEB;
		@(posedge clk8f);
		data_in_0 <= 'h26;
		data_in_1 <= 'hEA;
		@(posedge clk8f);
		data_in_0 <= 'h26;
		data_in_1 <= 'hEA;
		@(posedge clk8f);
		data_in_0 <= 'h26;
		data_in_1 <= 'hEA;
		@(posedge clk8f);
		data_in_0 <= 'h26;
		data_in_1 <= 'hEA;
		@(posedge clk8f);
		data_in_0 <= 'h26;
		data_in_1 <= 'hEA;
		@(posedge clk8f);
		data_in_0 <= 'h26;
		data_in_1 <= 'hEA;
		@(posedge clk8f);
		data_in_0 <= 'h26;
		data_in_1 <= 'hEA;
		@(posedge clk8f);
		data_in_0 <= 'h26;
		data_in_1 <= 'hEA;
		$finish;						// Termina de almacenar se�ales
	end
	// Reloj
	initial	clk8f 	<= 0;				// Valor inicial al reloj, sino siempre ser� indeterminado
	always	#45 clk8f 	<= ~clk8f;		// Hace "toggle" cada 2*10ns
	
endmodule
